module X ();

endmodule
