module X ();

endmodule
